library verilog;
use verilog.vl_types.all;
entity rgb_to_gray_vlg_vec_tst is
end rgb_to_gray_vlg_vec_tst;
